module sized_number_check;
